// megafunction wizard: %LPM_FIFO+%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: dcfifo 

// ============================================================
// File Name: Altera_UP_Video_In_Dual_Clock_FIFO.v
// Megafunction Name(s):
// 			dcfifo
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 6.1 Build 201 11/27/2006 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_up_video_dual_clock_fifo (
	// Inputs
	wrclk,
	wrreq,
	data,
	
	rdclk,
	rdreq,

	// Outputs	
	wrusedw,
	wrfull,

	q,
	rdusedw,
	rdempty
);

parameter DW = 18;

input				wrclk;
input				wrreq;
input	[(DW-1):0]  data;

input	 			rdclk;
input				rdreq;

output	[6:0]		wrusedw;
output				wrfull;

output	[(DW-1):0]	q;
output	[6:0]		rdusedw;
output				rdempty;

dcfifo	dcfifo_component (
	// Inputs
	.wrclk		(wrclk),
	.wrreq		(wrreq),
	.data		(data),
				
	.rdclk		(rdclk),
	.rdreq		(rdreq),

	// Outputs
	.wrusedw	(wrusedw),
	.wrfull		(wrfull),

	.q			(q),
	.rdusedw	(rdusedw),
	.rdempty	(rdempty)
	// synopsys translate_off
	,
	.aclr		(),
	.rdempty	(),
	.rdfull		(),
	.wrempty	()
	// synopsys translate_on
);
defparam
	dcfifo_component.intended_device_family	= "Cyclone II",
	dcfifo_component.lpm_hint				= "MAXIMIZE_SPEED=5,",
	dcfifo_component.lpm_numwords			= 128,
	dcfifo_component.lpm_showahead			= "ON",
	dcfifo_component.lpm_type				= "dcfifo",
	dcfifo_component.lpm_width				= DW,
	dcfifo_component.lpm_widthu				= 7,
	dcfifo_component.overflow_checking		= "ON",
	dcfifo_component.rdsync_delaypipe		= 4,
	dcfifo_component.underflow_checking		= "ON",
	dcfifo_component.use_eab				= "ON",
	dcfifo_component.wrsync_delaypipe		= 4;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AlmostEmpty NUMERIC "0"
// Retrieval info: PRIVATE: AlmostEmptyThr NUMERIC "-1"
// Retrieval info: PRIVATE: AlmostFull NUMERIC "0"
// Retrieval info: PRIVATE: AlmostFullThr NUMERIC "-1"
// Retrieval info: PRIVATE: CLOCKS_ARE_SYNCHRONIZED NUMERIC "0"
// Retrieval info: PRIVATE: Clock NUMERIC "4"
// Retrieval info: PRIVATE: Depth NUMERIC "128"
// Retrieval info: PRIVATE: Empty NUMERIC "1"
// Retrieval info: PRIVATE: Full NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: LE_BasedFIFO NUMERIC "0"
// Retrieval info: PRIVATE: LegacyRREQ NUMERIC "0"
// Retrieval info: PRIVATE: MAX_DEPTH_BY_9 NUMERIC "0"
// Retrieval info: PRIVATE: OVERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: Optimize NUMERIC "2"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: UNDERFLOW_CHECKING NUMERIC "0"
// Retrieval info: PRIVATE: UsedW NUMERIC "1"
// Retrieval info: PRIVATE: Width NUMERIC "26"
// Retrieval info: PRIVATE: dc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: diff_widths NUMERIC "0"
// Retrieval info: PRIVATE: output_width NUMERIC "26"
// Retrieval info: PRIVATE: rsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: rsFull NUMERIC "0"
// Retrieval info: PRIVATE: rsUsedW NUMERIC "1"
// Retrieval info: PRIVATE: sc_aclr NUMERIC "0"
// Retrieval info: PRIVATE: sc_sclr NUMERIC "0"
// Retrieval info: PRIVATE: wsEmpty NUMERIC "0"
// Retrieval info: PRIVATE: wsFull NUMERIC "0"
// Retrieval info: PRIVATE: wsUsedW NUMERIC "0"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=5,"
// Retrieval info: CONSTANT: LPM_NUMWORDS NUMERIC "128"
// Retrieval info: CONSTANT: LPM_SHOWAHEAD STRING "ON"
// Retrieval info: CONSTANT: LPM_TYPE STRING "dcfifo"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "26"
// Retrieval info: CONSTANT: LPM_WIDTHU NUMERIC "7"
// Retrieval info: CONSTANT: OVERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: RDSYNC_DELAYPIPE NUMERIC "4"
// Retrieval info: CONSTANT: UNDERFLOW_CHECKING STRING "ON"
// Retrieval info: CONSTANT: USE_EAB STRING "ON"
// Retrieval info: CONSTANT: WRSYNC_DELAYPIPE NUMERIC "4"
// Retrieval info: USED_PORT: data 0 0 26 0 INPUT NODEFVAL data[25..0]
// Retrieval info: USED_PORT: q 0 0 26 0 OUTPUT NODEFVAL q[25..0]
// Retrieval info: USED_PORT: rdclk 0 0 0 0 INPUT NODEFVAL rdclk
// Retrieval info: USED_PORT: rdreq 0 0 0 0 INPUT NODEFVAL rdreq
// Retrieval info: USED_PORT: rdusedw 0 0 7 0 OUTPUT NODEFVAL rdusedw[6..0]
// Retrieval info: USED_PORT: wrclk 0 0 0 0 INPUT NODEFVAL wrclk
// Retrieval info: USED_PORT: wrreq 0 0 0 0 INPUT NODEFVAL wrreq
// Retrieval info: CONNECT: @data 0 0 26 0 data 0 0 26 0
// Retrieval info: CONNECT: q 0 0 26 0 @q 0 0 26 0
// Retrieval info: CONNECT: @wrreq 0 0 0 0 wrreq 0 0 0 0
// Retrieval info: CONNECT: @rdreq 0 0 0 0 rdreq 0 0 0 0
// Retrieval info: CONNECT: @rdclk 0 0 0 0 rdclk 0 0 0 0
// Retrieval info: CONNECT: @wrclk 0 0 0 0 wrclk 0 0 0 0
// Retrieval info: CONNECT: rdusedw 0 0 7 0 @rdusedw 0 0 7 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL Altera_UP_Video_In_Dual_Clock_FIFO.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Altera_UP_Video_In_Dual_Clock_FIFO.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Altera_UP_Video_In_Dual_Clock_FIFO.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Altera_UP_Video_In_Dual_Clock_FIFO.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Altera_UP_Video_In_Dual_Clock_FIFO_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Altera_UP_Video_In_Dual_Clock_FIFO_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
